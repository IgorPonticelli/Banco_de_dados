-- Igor Ponticelli
-- igor.ponticelli@edu.pucrs.br

library ieee;
    use ieee.std_logic_1164.all;

entity somador_3b is
port
(
    op_a    :   in std_logic_vector(2 downto 0);
    op_b    :   in std_logic_vector(2 downto 0);
    soma    :   in std_logic_vector(3 downto 0)
);
end somador_3b;

architecture soma_maneira of somador_3b is

begin


end soma_maneira;